module mem_ext(
  input  [27:0] W0_addr,
  input         W0_clk,
  input  [63:0] W0_data,
  input         W0_en,
  input  [7:0]  W0_mask,
  input  [27:0] R0_addr,
  input         R0_clk,
  output [63:0] R0_data,
  input         R0_en
);
  wire [25:0] mem_0_0_W0_addr;
  wire  mem_0_0_W0_clk;
  wire [7:0] mem_0_0_W0_data;
  wire  mem_0_0_W0_en;
  wire  mem_0_0_W0_mask;
  wire [25:0] mem_0_0_R0_addr;
  wire  mem_0_0_R0_clk;
  wire [7:0] mem_0_0_R0_data;
  wire  mem_0_0_R0_en;
  wire [25:0] mem_0_1_W0_addr;
  wire  mem_0_1_W0_clk;
  wire [7:0] mem_0_1_W0_data;
  wire  mem_0_1_W0_en;
  wire  mem_0_1_W0_mask;
  wire [25:0] mem_0_1_R0_addr;
  wire  mem_0_1_R0_clk;
  wire [7:0] mem_0_1_R0_data;
  wire  mem_0_1_R0_en;
  wire [25:0] mem_0_2_W0_addr;
  wire  mem_0_2_W0_clk;
  wire [7:0] mem_0_2_W0_data;
  wire  mem_0_2_W0_en;
  wire  mem_0_2_W0_mask;
  wire [25:0] mem_0_2_R0_addr;
  wire  mem_0_2_R0_clk;
  wire [7:0] mem_0_2_R0_data;
  wire  mem_0_2_R0_en;
  wire [25:0] mem_0_3_W0_addr;
  wire  mem_0_3_W0_clk;
  wire [7:0] mem_0_3_W0_data;
  wire  mem_0_3_W0_en;
  wire  mem_0_3_W0_mask;
  wire [25:0] mem_0_3_R0_addr;
  wire  mem_0_3_R0_clk;
  wire [7:0] mem_0_3_R0_data;
  wire  mem_0_3_R0_en;
  wire [25:0] mem_0_4_W0_addr;
  wire  mem_0_4_W0_clk;
  wire [7:0] mem_0_4_W0_data;
  wire  mem_0_4_W0_en;
  wire  mem_0_4_W0_mask;
  wire [25:0] mem_0_4_R0_addr;
  wire  mem_0_4_R0_clk;
  wire [7:0] mem_0_4_R0_data;
  wire  mem_0_4_R0_en;
  wire [25:0] mem_0_5_W0_addr;
  wire  mem_0_5_W0_clk;
  wire [7:0] mem_0_5_W0_data;
  wire  mem_0_5_W0_en;
  wire  mem_0_5_W0_mask;
  wire [25:0] mem_0_5_R0_addr;
  wire  mem_0_5_R0_clk;
  wire [7:0] mem_0_5_R0_data;
  wire  mem_0_5_R0_en;
  wire [25:0] mem_0_6_W0_addr;
  wire  mem_0_6_W0_clk;
  wire [7:0] mem_0_6_W0_data;
  wire  mem_0_6_W0_en;
  wire  mem_0_6_W0_mask;
  wire [25:0] mem_0_6_R0_addr;
  wire  mem_0_6_R0_clk;
  wire [7:0] mem_0_6_R0_data;
  wire  mem_0_6_R0_en;
  wire [25:0] mem_0_7_W0_addr;
  wire  mem_0_7_W0_clk;
  wire [7:0] mem_0_7_W0_data;
  wire  mem_0_7_W0_en;
  wire  mem_0_7_W0_mask;
  wire [25:0] mem_0_7_R0_addr;
  wire  mem_0_7_R0_clk;
  wire [7:0] mem_0_7_R0_data;
  wire  mem_0_7_R0_en;
  wire [25:0] mem_1_0_W0_addr;
  wire  mem_1_0_W0_clk;
  wire [7:0] mem_1_0_W0_data;
  wire  mem_1_0_W0_en;
  wire  mem_1_0_W0_mask;
  wire [25:0] mem_1_0_R0_addr;
  wire  mem_1_0_R0_clk;
  wire [7:0] mem_1_0_R0_data;
  wire  mem_1_0_R0_en;
  wire [25:0] mem_1_1_W0_addr;
  wire  mem_1_1_W0_clk;
  wire [7:0] mem_1_1_W0_data;
  wire  mem_1_1_W0_en;
  wire  mem_1_1_W0_mask;
  wire [25:0] mem_1_1_R0_addr;
  wire  mem_1_1_R0_clk;
  wire [7:0] mem_1_1_R0_data;
  wire  mem_1_1_R0_en;
  wire [25:0] mem_1_2_W0_addr;
  wire  mem_1_2_W0_clk;
  wire [7:0] mem_1_2_W0_data;
  wire  mem_1_2_W0_en;
  wire  mem_1_2_W0_mask;
  wire [25:0] mem_1_2_R0_addr;
  wire  mem_1_2_R0_clk;
  wire [7:0] mem_1_2_R0_data;
  wire  mem_1_2_R0_en;
  wire [25:0] mem_1_3_W0_addr;
  wire  mem_1_3_W0_clk;
  wire [7:0] mem_1_3_W0_data;
  wire  mem_1_3_W0_en;
  wire  mem_1_3_W0_mask;
  wire [25:0] mem_1_3_R0_addr;
  wire  mem_1_3_R0_clk;
  wire [7:0] mem_1_3_R0_data;
  wire  mem_1_3_R0_en;
  wire [25:0] mem_1_4_W0_addr;
  wire  mem_1_4_W0_clk;
  wire [7:0] mem_1_4_W0_data;
  wire  mem_1_4_W0_en;
  wire  mem_1_4_W0_mask;
  wire [25:0] mem_1_4_R0_addr;
  wire  mem_1_4_R0_clk;
  wire [7:0] mem_1_4_R0_data;
  wire  mem_1_4_R0_en;
  wire [25:0] mem_1_5_W0_addr;
  wire  mem_1_5_W0_clk;
  wire [7:0] mem_1_5_W0_data;
  wire  mem_1_5_W0_en;
  wire  mem_1_5_W0_mask;
  wire [25:0] mem_1_5_R0_addr;
  wire  mem_1_5_R0_clk;
  wire [7:0] mem_1_5_R0_data;
  wire  mem_1_5_R0_en;
  wire [25:0] mem_1_6_W0_addr;
  wire  mem_1_6_W0_clk;
  wire [7:0] mem_1_6_W0_data;
  wire  mem_1_6_W0_en;
  wire  mem_1_6_W0_mask;
  wire [25:0] mem_1_6_R0_addr;
  wire  mem_1_6_R0_clk;
  wire [7:0] mem_1_6_R0_data;
  wire  mem_1_6_R0_en;
  wire [25:0] mem_1_7_W0_addr;
  wire  mem_1_7_W0_clk;
  wire [7:0] mem_1_7_W0_data;
  wire  mem_1_7_W0_en;
  wire  mem_1_7_W0_mask;
  wire [25:0] mem_1_7_R0_addr;
  wire  mem_1_7_R0_clk;
  wire [7:0] mem_1_7_R0_data;
  wire  mem_1_7_R0_en;
  wire [25:0] mem_2_0_W0_addr;
  wire  mem_2_0_W0_clk;
  wire [7:0] mem_2_0_W0_data;
  wire  mem_2_0_W0_en;
  wire  mem_2_0_W0_mask;
  wire [25:0] mem_2_0_R0_addr;
  wire  mem_2_0_R0_clk;
  wire [7:0] mem_2_0_R0_data;
  wire  mem_2_0_R0_en;
  wire [25:0] mem_2_1_W0_addr;
  wire  mem_2_1_W0_clk;
  wire [7:0] mem_2_1_W0_data;
  wire  mem_2_1_W0_en;
  wire  mem_2_1_W0_mask;
  wire [25:0] mem_2_1_R0_addr;
  wire  mem_2_1_R0_clk;
  wire [7:0] mem_2_1_R0_data;
  wire  mem_2_1_R0_en;
  wire [25:0] mem_2_2_W0_addr;
  wire  mem_2_2_W0_clk;
  wire [7:0] mem_2_2_W0_data;
  wire  mem_2_2_W0_en;
  wire  mem_2_2_W0_mask;
  wire [25:0] mem_2_2_R0_addr;
  wire  mem_2_2_R0_clk;
  wire [7:0] mem_2_2_R0_data;
  wire  mem_2_2_R0_en;
  wire [25:0] mem_2_3_W0_addr;
  wire  mem_2_3_W0_clk;
  wire [7:0] mem_2_3_W0_data;
  wire  mem_2_3_W0_en;
  wire  mem_2_3_W0_mask;
  wire [25:0] mem_2_3_R0_addr;
  wire  mem_2_3_R0_clk;
  wire [7:0] mem_2_3_R0_data;
  wire  mem_2_3_R0_en;
  wire [25:0] mem_2_4_W0_addr;
  wire  mem_2_4_W0_clk;
  wire [7:0] mem_2_4_W0_data;
  wire  mem_2_4_W0_en;
  wire  mem_2_4_W0_mask;
  wire [25:0] mem_2_4_R0_addr;
  wire  mem_2_4_R0_clk;
  wire [7:0] mem_2_4_R0_data;
  wire  mem_2_4_R0_en;
  wire [25:0] mem_2_5_W0_addr;
  wire  mem_2_5_W0_clk;
  wire [7:0] mem_2_5_W0_data;
  wire  mem_2_5_W0_en;
  wire  mem_2_5_W0_mask;
  wire [25:0] mem_2_5_R0_addr;
  wire  mem_2_5_R0_clk;
  wire [7:0] mem_2_5_R0_data;
  wire  mem_2_5_R0_en;
  wire [25:0] mem_2_6_W0_addr;
  wire  mem_2_6_W0_clk;
  wire [7:0] mem_2_6_W0_data;
  wire  mem_2_6_W0_en;
  wire  mem_2_6_W0_mask;
  wire [25:0] mem_2_6_R0_addr;
  wire  mem_2_6_R0_clk;
  wire [7:0] mem_2_6_R0_data;
  wire  mem_2_6_R0_en;
  wire [25:0] mem_2_7_W0_addr;
  wire  mem_2_7_W0_clk;
  wire [7:0] mem_2_7_W0_data;
  wire  mem_2_7_W0_en;
  wire  mem_2_7_W0_mask;
  wire [25:0] mem_2_7_R0_addr;
  wire  mem_2_7_R0_clk;
  wire [7:0] mem_2_7_R0_data;
  wire  mem_2_7_R0_en;
  wire [25:0] mem_3_0_W0_addr;
  wire  mem_3_0_W0_clk;
  wire [7:0] mem_3_0_W0_data;
  wire  mem_3_0_W0_en;
  wire  mem_3_0_W0_mask;
  wire [25:0] mem_3_0_R0_addr;
  wire  mem_3_0_R0_clk;
  wire [7:0] mem_3_0_R0_data;
  wire  mem_3_0_R0_en;
  wire [25:0] mem_3_1_W0_addr;
  wire  mem_3_1_W0_clk;
  wire [7:0] mem_3_1_W0_data;
  wire  mem_3_1_W0_en;
  wire  mem_3_1_W0_mask;
  wire [25:0] mem_3_1_R0_addr;
  wire  mem_3_1_R0_clk;
  wire [7:0] mem_3_1_R0_data;
  wire  mem_3_1_R0_en;
  wire [25:0] mem_3_2_W0_addr;
  wire  mem_3_2_W0_clk;
  wire [7:0] mem_3_2_W0_data;
  wire  mem_3_2_W0_en;
  wire  mem_3_2_W0_mask;
  wire [25:0] mem_3_2_R0_addr;
  wire  mem_3_2_R0_clk;
  wire [7:0] mem_3_2_R0_data;
  wire  mem_3_2_R0_en;
  wire [25:0] mem_3_3_W0_addr;
  wire  mem_3_3_W0_clk;
  wire [7:0] mem_3_3_W0_data;
  wire  mem_3_3_W0_en;
  wire  mem_3_3_W0_mask;
  wire [25:0] mem_3_3_R0_addr;
  wire  mem_3_3_R0_clk;
  wire [7:0] mem_3_3_R0_data;
  wire  mem_3_3_R0_en;
  wire [25:0] mem_3_4_W0_addr;
  wire  mem_3_4_W0_clk;
  wire [7:0] mem_3_4_W0_data;
  wire  mem_3_4_W0_en;
  wire  mem_3_4_W0_mask;
  wire [25:0] mem_3_4_R0_addr;
  wire  mem_3_4_R0_clk;
  wire [7:0] mem_3_4_R0_data;
  wire  mem_3_4_R0_en;
  wire [25:0] mem_3_5_W0_addr;
  wire  mem_3_5_W0_clk;
  wire [7:0] mem_3_5_W0_data;
  wire  mem_3_5_W0_en;
  wire  mem_3_5_W0_mask;
  wire [25:0] mem_3_5_R0_addr;
  wire  mem_3_5_R0_clk;
  wire [7:0] mem_3_5_R0_data;
  wire  mem_3_5_R0_en;
  wire [25:0] mem_3_6_W0_addr;
  wire  mem_3_6_W0_clk;
  wire [7:0] mem_3_6_W0_data;
  wire  mem_3_6_W0_en;
  wire  mem_3_6_W0_mask;
  wire [25:0] mem_3_6_R0_addr;
  wire  mem_3_6_R0_clk;
  wire [7:0] mem_3_6_R0_data;
  wire  mem_3_6_R0_en;
  wire [25:0] mem_3_7_W0_addr;
  wire  mem_3_7_W0_clk;
  wire [7:0] mem_3_7_W0_data;
  wire  mem_3_7_W0_en;
  wire  mem_3_7_W0_mask;
  wire [25:0] mem_3_7_R0_addr;
  wire  mem_3_7_R0_clk;
  wire [7:0] mem_3_7_R0_data;
  wire  mem_3_7_R0_en;
  wire [1:0] W0_addr_sel;
  wire [1:0] R0_addr_sel;
  reg [1:0] R0_addr_sel_reg;
  reg [31:0] _RAND_0;
  wire [7:0] R0_data_0_0;
  wire [7:0] R0_data_0_1;
  wire [7:0] R0_data_0_2;
  wire [7:0] R0_data_0_3;
  wire [7:0] R0_data_0_4;
  wire [7:0] R0_data_0_5;
  wire [7:0] R0_data_0_6;
  wire [7:0] R0_data_0_7;
  wire [15:0] _GEN_0;
  wire [23:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire [39:0] _GEN_3;
  wire [47:0] _GEN_4;
  wire [55:0] _GEN_5;
  wire [63:0] R0_data_0;
  wire [7:0] R0_data_1_0;
  wire [7:0] R0_data_1_1;
  wire [7:0] R0_data_1_2;
  wire [7:0] R0_data_1_3;
  wire [7:0] R0_data_1_4;
  wire [7:0] R0_data_1_5;
  wire [7:0] R0_data_1_6;
  wire [7:0] R0_data_1_7;
  wire [15:0] _GEN_6;
  wire [23:0] _GEN_7;
  wire [31:0] _GEN_8;
  wire [39:0] _GEN_9;
  wire [47:0] _GEN_10;
  wire [55:0] _GEN_11;
  wire [63:0] R0_data_1;
  wire [7:0] R0_data_2_0;
  wire [7:0] R0_data_2_1;
  wire [7:0] R0_data_2_2;
  wire [7:0] R0_data_2_3;
  wire [7:0] R0_data_2_4;
  wire [7:0] R0_data_2_5;
  wire [7:0] R0_data_2_6;
  wire [7:0] R0_data_2_7;
  wire [15:0] _GEN_12;
  wire [23:0] _GEN_13;
  wire [31:0] _GEN_14;
  wire [39:0] _GEN_15;
  wire [47:0] _GEN_16;
  wire [55:0] _GEN_17;
  wire [63:0] R0_data_2;
  wire [7:0] R0_data_3_0;
  wire [7:0] R0_data_3_1;
  wire [7:0] R0_data_3_2;
  wire [7:0] R0_data_3_3;
  wire [7:0] R0_data_3_4;
  wire [7:0] R0_data_3_5;
  wire [7:0] R0_data_3_6;
  wire [7:0] R0_data_3_7;
  wire [15:0] _GEN_18;
  wire [23:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire [39:0] _GEN_21;
  wire [47:0] _GEN_22;
  wire [55:0] _GEN_23;
  wire [63:0] R0_data_3;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire  _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_76;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire  _GEN_83;
  wire  _GEN_84;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _GEN_87;
  split_mem_ext mem_0_0 (
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_mem_ext mem_0_1 (
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_mem_ext mem_0_2 (
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_mem_ext mem_0_3 (
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  split_mem_ext mem_0_4 (
    .W0_addr(mem_0_4_W0_addr),
    .W0_clk(mem_0_4_W0_clk),
    .W0_data(mem_0_4_W0_data),
    .W0_en(mem_0_4_W0_en),
    .W0_mask(mem_0_4_W0_mask),
    .R0_addr(mem_0_4_R0_addr),
    .R0_clk(mem_0_4_R0_clk),
    .R0_data(mem_0_4_R0_data),
    .R0_en(mem_0_4_R0_en)
  );
  split_mem_ext mem_0_5 (
    .W0_addr(mem_0_5_W0_addr),
    .W0_clk(mem_0_5_W0_clk),
    .W0_data(mem_0_5_W0_data),
    .W0_en(mem_0_5_W0_en),
    .W0_mask(mem_0_5_W0_mask),
    .R0_addr(mem_0_5_R0_addr),
    .R0_clk(mem_0_5_R0_clk),
    .R0_data(mem_0_5_R0_data),
    .R0_en(mem_0_5_R0_en)
  );
  split_mem_ext mem_0_6 (
    .W0_addr(mem_0_6_W0_addr),
    .W0_clk(mem_0_6_W0_clk),
    .W0_data(mem_0_6_W0_data),
    .W0_en(mem_0_6_W0_en),
    .W0_mask(mem_0_6_W0_mask),
    .R0_addr(mem_0_6_R0_addr),
    .R0_clk(mem_0_6_R0_clk),
    .R0_data(mem_0_6_R0_data),
    .R0_en(mem_0_6_R0_en)
  );
  split_mem_ext mem_0_7 (
    .W0_addr(mem_0_7_W0_addr),
    .W0_clk(mem_0_7_W0_clk),
    .W0_data(mem_0_7_W0_data),
    .W0_en(mem_0_7_W0_en),
    .W0_mask(mem_0_7_W0_mask),
    .R0_addr(mem_0_7_R0_addr),
    .R0_clk(mem_0_7_R0_clk),
    .R0_data(mem_0_7_R0_data),
    .R0_en(mem_0_7_R0_en)
  );
  split_mem_ext mem_1_0 (
    .W0_addr(mem_1_0_W0_addr),
    .W0_clk(mem_1_0_W0_clk),
    .W0_data(mem_1_0_W0_data),
    .W0_en(mem_1_0_W0_en),
    .W0_mask(mem_1_0_W0_mask),
    .R0_addr(mem_1_0_R0_addr),
    .R0_clk(mem_1_0_R0_clk),
    .R0_data(mem_1_0_R0_data),
    .R0_en(mem_1_0_R0_en)
  );
  split_mem_ext mem_1_1 (
    .W0_addr(mem_1_1_W0_addr),
    .W0_clk(mem_1_1_W0_clk),
    .W0_data(mem_1_1_W0_data),
    .W0_en(mem_1_1_W0_en),
    .W0_mask(mem_1_1_W0_mask),
    .R0_addr(mem_1_1_R0_addr),
    .R0_clk(mem_1_1_R0_clk),
    .R0_data(mem_1_1_R0_data),
    .R0_en(mem_1_1_R0_en)
  );
  split_mem_ext mem_1_2 (
    .W0_addr(mem_1_2_W0_addr),
    .W0_clk(mem_1_2_W0_clk),
    .W0_data(mem_1_2_W0_data),
    .W0_en(mem_1_2_W0_en),
    .W0_mask(mem_1_2_W0_mask),
    .R0_addr(mem_1_2_R0_addr),
    .R0_clk(mem_1_2_R0_clk),
    .R0_data(mem_1_2_R0_data),
    .R0_en(mem_1_2_R0_en)
  );
  split_mem_ext mem_1_3 (
    .W0_addr(mem_1_3_W0_addr),
    .W0_clk(mem_1_3_W0_clk),
    .W0_data(mem_1_3_W0_data),
    .W0_en(mem_1_3_W0_en),
    .W0_mask(mem_1_3_W0_mask),
    .R0_addr(mem_1_3_R0_addr),
    .R0_clk(mem_1_3_R0_clk),
    .R0_data(mem_1_3_R0_data),
    .R0_en(mem_1_3_R0_en)
  );
  split_mem_ext mem_1_4 (
    .W0_addr(mem_1_4_W0_addr),
    .W0_clk(mem_1_4_W0_clk),
    .W0_data(mem_1_4_W0_data),
    .W0_en(mem_1_4_W0_en),
    .W0_mask(mem_1_4_W0_mask),
    .R0_addr(mem_1_4_R0_addr),
    .R0_clk(mem_1_4_R0_clk),
    .R0_data(mem_1_4_R0_data),
    .R0_en(mem_1_4_R0_en)
  );
  split_mem_ext mem_1_5 (
    .W0_addr(mem_1_5_W0_addr),
    .W0_clk(mem_1_5_W0_clk),
    .W0_data(mem_1_5_W0_data),
    .W0_en(mem_1_5_W0_en),
    .W0_mask(mem_1_5_W0_mask),
    .R0_addr(mem_1_5_R0_addr),
    .R0_clk(mem_1_5_R0_clk),
    .R0_data(mem_1_5_R0_data),
    .R0_en(mem_1_5_R0_en)
  );
  split_mem_ext mem_1_6 (
    .W0_addr(mem_1_6_W0_addr),
    .W0_clk(mem_1_6_W0_clk),
    .W0_data(mem_1_6_W0_data),
    .W0_en(mem_1_6_W0_en),
    .W0_mask(mem_1_6_W0_mask),
    .R0_addr(mem_1_6_R0_addr),
    .R0_clk(mem_1_6_R0_clk),
    .R0_data(mem_1_6_R0_data),
    .R0_en(mem_1_6_R0_en)
  );
  split_mem_ext mem_1_7 (
    .W0_addr(mem_1_7_W0_addr),
    .W0_clk(mem_1_7_W0_clk),
    .W0_data(mem_1_7_W0_data),
    .W0_en(mem_1_7_W0_en),
    .W0_mask(mem_1_7_W0_mask),
    .R0_addr(mem_1_7_R0_addr),
    .R0_clk(mem_1_7_R0_clk),
    .R0_data(mem_1_7_R0_data),
    .R0_en(mem_1_7_R0_en)
  );
  split_mem_ext mem_2_0 (
    .W0_addr(mem_2_0_W0_addr),
    .W0_clk(mem_2_0_W0_clk),
    .W0_data(mem_2_0_W0_data),
    .W0_en(mem_2_0_W0_en),
    .W0_mask(mem_2_0_W0_mask),
    .R0_addr(mem_2_0_R0_addr),
    .R0_clk(mem_2_0_R0_clk),
    .R0_data(mem_2_0_R0_data),
    .R0_en(mem_2_0_R0_en)
  );
  split_mem_ext mem_2_1 (
    .W0_addr(mem_2_1_W0_addr),
    .W0_clk(mem_2_1_W0_clk),
    .W0_data(mem_2_1_W0_data),
    .W0_en(mem_2_1_W0_en),
    .W0_mask(mem_2_1_W0_mask),
    .R0_addr(mem_2_1_R0_addr),
    .R0_clk(mem_2_1_R0_clk),
    .R0_data(mem_2_1_R0_data),
    .R0_en(mem_2_1_R0_en)
  );
  split_mem_ext mem_2_2 (
    .W0_addr(mem_2_2_W0_addr),
    .W0_clk(mem_2_2_W0_clk),
    .W0_data(mem_2_2_W0_data),
    .W0_en(mem_2_2_W0_en),
    .W0_mask(mem_2_2_W0_mask),
    .R0_addr(mem_2_2_R0_addr),
    .R0_clk(mem_2_2_R0_clk),
    .R0_data(mem_2_2_R0_data),
    .R0_en(mem_2_2_R0_en)
  );
  split_mem_ext mem_2_3 (
    .W0_addr(mem_2_3_W0_addr),
    .W0_clk(mem_2_3_W0_clk),
    .W0_data(mem_2_3_W0_data),
    .W0_en(mem_2_3_W0_en),
    .W0_mask(mem_2_3_W0_mask),
    .R0_addr(mem_2_3_R0_addr),
    .R0_clk(mem_2_3_R0_clk),
    .R0_data(mem_2_3_R0_data),
    .R0_en(mem_2_3_R0_en)
  );
  split_mem_ext mem_2_4 (
    .W0_addr(mem_2_4_W0_addr),
    .W0_clk(mem_2_4_W0_clk),
    .W0_data(mem_2_4_W0_data),
    .W0_en(mem_2_4_W0_en),
    .W0_mask(mem_2_4_W0_mask),
    .R0_addr(mem_2_4_R0_addr),
    .R0_clk(mem_2_4_R0_clk),
    .R0_data(mem_2_4_R0_data),
    .R0_en(mem_2_4_R0_en)
  );
  split_mem_ext mem_2_5 (
    .W0_addr(mem_2_5_W0_addr),
    .W0_clk(mem_2_5_W0_clk),
    .W0_data(mem_2_5_W0_data),
    .W0_en(mem_2_5_W0_en),
    .W0_mask(mem_2_5_W0_mask),
    .R0_addr(mem_2_5_R0_addr),
    .R0_clk(mem_2_5_R0_clk),
    .R0_data(mem_2_5_R0_data),
    .R0_en(mem_2_5_R0_en)
  );
  split_mem_ext mem_2_6 (
    .W0_addr(mem_2_6_W0_addr),
    .W0_clk(mem_2_6_W0_clk),
    .W0_data(mem_2_6_W0_data),
    .W0_en(mem_2_6_W0_en),
    .W0_mask(mem_2_6_W0_mask),
    .R0_addr(mem_2_6_R0_addr),
    .R0_clk(mem_2_6_R0_clk),
    .R0_data(mem_2_6_R0_data),
    .R0_en(mem_2_6_R0_en)
  );
  split_mem_ext mem_2_7 (
    .W0_addr(mem_2_7_W0_addr),
    .W0_clk(mem_2_7_W0_clk),
    .W0_data(mem_2_7_W0_data),
    .W0_en(mem_2_7_W0_en),
    .W0_mask(mem_2_7_W0_mask),
    .R0_addr(mem_2_7_R0_addr),
    .R0_clk(mem_2_7_R0_clk),
    .R0_data(mem_2_7_R0_data),
    .R0_en(mem_2_7_R0_en)
  );
  split_mem_ext mem_3_0 (
    .W0_addr(mem_3_0_W0_addr),
    .W0_clk(mem_3_0_W0_clk),
    .W0_data(mem_3_0_W0_data),
    .W0_en(mem_3_0_W0_en),
    .W0_mask(mem_3_0_W0_mask),
    .R0_addr(mem_3_0_R0_addr),
    .R0_clk(mem_3_0_R0_clk),
    .R0_data(mem_3_0_R0_data),
    .R0_en(mem_3_0_R0_en)
  );
  split_mem_ext mem_3_1 (
    .W0_addr(mem_3_1_W0_addr),
    .W0_clk(mem_3_1_W0_clk),
    .W0_data(mem_3_1_W0_data),
    .W0_en(mem_3_1_W0_en),
    .W0_mask(mem_3_1_W0_mask),
    .R0_addr(mem_3_1_R0_addr),
    .R0_clk(mem_3_1_R0_clk),
    .R0_data(mem_3_1_R0_data),
    .R0_en(mem_3_1_R0_en)
  );
  split_mem_ext mem_3_2 (
    .W0_addr(mem_3_2_W0_addr),
    .W0_clk(mem_3_2_W0_clk),
    .W0_data(mem_3_2_W0_data),
    .W0_en(mem_3_2_W0_en),
    .W0_mask(mem_3_2_W0_mask),
    .R0_addr(mem_3_2_R0_addr),
    .R0_clk(mem_3_2_R0_clk),
    .R0_data(mem_3_2_R0_data),
    .R0_en(mem_3_2_R0_en)
  );
  split_mem_ext mem_3_3 (
    .W0_addr(mem_3_3_W0_addr),
    .W0_clk(mem_3_3_W0_clk),
    .W0_data(mem_3_3_W0_data),
    .W0_en(mem_3_3_W0_en),
    .W0_mask(mem_3_3_W0_mask),
    .R0_addr(mem_3_3_R0_addr),
    .R0_clk(mem_3_3_R0_clk),
    .R0_data(mem_3_3_R0_data),
    .R0_en(mem_3_3_R0_en)
  );
  split_mem_ext mem_3_4 (
    .W0_addr(mem_3_4_W0_addr),
    .W0_clk(mem_3_4_W0_clk),
    .W0_data(mem_3_4_W0_data),
    .W0_en(mem_3_4_W0_en),
    .W0_mask(mem_3_4_W0_mask),
    .R0_addr(mem_3_4_R0_addr),
    .R0_clk(mem_3_4_R0_clk),
    .R0_data(mem_3_4_R0_data),
    .R0_en(mem_3_4_R0_en)
  );
  split_mem_ext mem_3_5 (
    .W0_addr(mem_3_5_W0_addr),
    .W0_clk(mem_3_5_W0_clk),
    .W0_data(mem_3_5_W0_data),
    .W0_en(mem_3_5_W0_en),
    .W0_mask(mem_3_5_W0_mask),
    .R0_addr(mem_3_5_R0_addr),
    .R0_clk(mem_3_5_R0_clk),
    .R0_data(mem_3_5_R0_data),
    .R0_en(mem_3_5_R0_en)
  );
  split_mem_ext mem_3_6 (
    .W0_addr(mem_3_6_W0_addr),
    .W0_clk(mem_3_6_W0_clk),
    .W0_data(mem_3_6_W0_data),
    .W0_en(mem_3_6_W0_en),
    .W0_mask(mem_3_6_W0_mask),
    .R0_addr(mem_3_6_R0_addr),
    .R0_clk(mem_3_6_R0_clk),
    .R0_data(mem_3_6_R0_data),
    .R0_en(mem_3_6_R0_en)
  );
  split_mem_ext mem_3_7 (
    .W0_addr(mem_3_7_W0_addr),
    .W0_clk(mem_3_7_W0_clk),
    .W0_data(mem_3_7_W0_data),
    .W0_en(mem_3_7_W0_en),
    .W0_mask(mem_3_7_W0_mask),
    .R0_addr(mem_3_7_R0_addr),
    .R0_clk(mem_3_7_R0_clk),
    .R0_data(mem_3_7_R0_data),
    .R0_en(mem_3_7_R0_en)
  );
  assign W0_addr_sel = W0_addr[27:26];
  assign R0_addr_sel = R0_addr[27:26];
  assign R0_data_0_0 = mem_0_0_R0_data;
  assign R0_data_0_1 = mem_0_1_R0_data;
  assign R0_data_0_2 = mem_0_2_R0_data;
  assign R0_data_0_3 = mem_0_3_R0_data;
  assign R0_data_0_4 = mem_0_4_R0_data;
  assign R0_data_0_5 = mem_0_5_R0_data;
  assign R0_data_0_6 = mem_0_6_R0_data;
  assign R0_data_0_7 = mem_0_7_R0_data;
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0};
  assign _GEN_1 = {R0_data_0_2,_GEN_0};
  assign _GEN_2 = {R0_data_0_3,_GEN_1};
  assign _GEN_3 = {R0_data_0_4,_GEN_2};
  assign _GEN_4 = {R0_data_0_5,_GEN_3};
  assign _GEN_5 = {R0_data_0_6,_GEN_4};
  assign R0_data_0 = {R0_data_0_7,_GEN_5};
  assign R0_data_1_0 = mem_1_0_R0_data;
  assign R0_data_1_1 = mem_1_1_R0_data;
  assign R0_data_1_2 = mem_1_2_R0_data;
  assign R0_data_1_3 = mem_1_3_R0_data;
  assign R0_data_1_4 = mem_1_4_R0_data;
  assign R0_data_1_5 = mem_1_5_R0_data;
  assign R0_data_1_6 = mem_1_6_R0_data;
  assign R0_data_1_7 = mem_1_7_R0_data;
  assign _GEN_6 = {R0_data_1_1,R0_data_1_0};
  assign _GEN_7 = {R0_data_1_2,_GEN_6};
  assign _GEN_8 = {R0_data_1_3,_GEN_7};
  assign _GEN_9 = {R0_data_1_4,_GEN_8};
  assign _GEN_10 = {R0_data_1_5,_GEN_9};
  assign _GEN_11 = {R0_data_1_6,_GEN_10};
  assign R0_data_1 = {R0_data_1_7,_GEN_11};
  assign R0_data_2_0 = mem_2_0_R0_data;
  assign R0_data_2_1 = mem_2_1_R0_data;
  assign R0_data_2_2 = mem_2_2_R0_data;
  assign R0_data_2_3 = mem_2_3_R0_data;
  assign R0_data_2_4 = mem_2_4_R0_data;
  assign R0_data_2_5 = mem_2_5_R0_data;
  assign R0_data_2_6 = mem_2_6_R0_data;
  assign R0_data_2_7 = mem_2_7_R0_data;
  assign _GEN_12 = {R0_data_2_1,R0_data_2_0};
  assign _GEN_13 = {R0_data_2_2,_GEN_12};
  assign _GEN_14 = {R0_data_2_3,_GEN_13};
  assign _GEN_15 = {R0_data_2_4,_GEN_14};
  assign _GEN_16 = {R0_data_2_5,_GEN_15};
  assign _GEN_17 = {R0_data_2_6,_GEN_16};
  assign R0_data_2 = {R0_data_2_7,_GEN_17};
  assign R0_data_3_0 = mem_3_0_R0_data;
  assign R0_data_3_1 = mem_3_1_R0_data;
  assign R0_data_3_2 = mem_3_2_R0_data;
  assign R0_data_3_3 = mem_3_3_R0_data;
  assign R0_data_3_4 = mem_3_4_R0_data;
  assign R0_data_3_5 = mem_3_5_R0_data;
  assign R0_data_3_6 = mem_3_6_R0_data;
  assign R0_data_3_7 = mem_3_7_R0_data;
  assign _GEN_18 = {R0_data_3_1,R0_data_3_0};
  assign _GEN_19 = {R0_data_3_2,_GEN_18};
  assign _GEN_20 = {R0_data_3_3,_GEN_19};
  assign _GEN_21 = {R0_data_3_4,_GEN_20};
  assign _GEN_22 = {R0_data_3_5,_GEN_21};
  assign _GEN_23 = {R0_data_3_6,_GEN_22};
  assign R0_data_3 = {R0_data_3_7,_GEN_23};
  assign R0_data = R0_addr_sel_reg == 2'h0 ? R0_data_0 : R0_addr_sel_reg == 2'h1 ? R0_data_1 : R0_addr_sel_reg == 2'h2 ? R0_data_2 : R0_addr_sel_reg == 2'h3 ? R0_data_3 : 1'h0;
  assign mem_0_0_W0_addr = W0_addr[25:0];
  assign mem_0_0_W0_clk = W0_clk;
  assign mem_0_0_W0_data = W0_data[7:0];
  assign _GEN_24 = W0_addr_sel == 2'h0;
  assign mem_0_0_W0_en = W0_en & _GEN_24;
  assign mem_0_0_W0_mask = W0_mask[0];
  assign mem_0_0_R0_addr = R0_addr[25:0];
  assign mem_0_0_R0_clk = R0_clk;
  assign _GEN_25 = R0_addr_sel == 2'h0;
  assign mem_0_0_R0_en = R0_en & _GEN_25;
  assign mem_0_1_W0_addr = W0_addr[25:0];
  assign mem_0_1_W0_clk = W0_clk;
  assign mem_0_1_W0_data = W0_data[15:8];
  assign _GEN_26 = W0_addr_sel == 2'h0;
  assign mem_0_1_W0_en = W0_en & _GEN_24;
  assign mem_0_1_W0_mask = W0_mask[1];
  assign mem_0_1_R0_addr = R0_addr[25:0];
  assign mem_0_1_R0_clk = R0_clk;
  assign _GEN_27 = R0_addr_sel == 2'h0;
  assign mem_0_1_R0_en = R0_en & _GEN_25;
  assign mem_0_2_W0_addr = W0_addr[25:0];
  assign mem_0_2_W0_clk = W0_clk;
  assign mem_0_2_W0_data = W0_data[23:16];
  assign _GEN_28 = W0_addr_sel == 2'h0;
  assign mem_0_2_W0_en = W0_en & _GEN_24;
  assign mem_0_2_W0_mask = W0_mask[2];
  assign mem_0_2_R0_addr = R0_addr[25:0];
  assign mem_0_2_R0_clk = R0_clk;
  assign _GEN_29 = R0_addr_sel == 2'h0;
  assign mem_0_2_R0_en = R0_en & _GEN_25;
  assign mem_0_3_W0_addr = W0_addr[25:0];
  assign mem_0_3_W0_clk = W0_clk;
  assign mem_0_3_W0_data = W0_data[31:24];
  assign _GEN_30 = W0_addr_sel == 2'h0;
  assign mem_0_3_W0_en = W0_en & _GEN_24;
  assign mem_0_3_W0_mask = W0_mask[3];
  assign mem_0_3_R0_addr = R0_addr[25:0];
  assign mem_0_3_R0_clk = R0_clk;
  assign _GEN_31 = R0_addr_sel == 2'h0;
  assign mem_0_3_R0_en = R0_en & _GEN_25;
  assign mem_0_4_W0_addr = W0_addr[25:0];
  assign mem_0_4_W0_clk = W0_clk;
  assign mem_0_4_W0_data = W0_data[39:32];
  assign _GEN_32 = W0_addr_sel == 2'h0;
  assign mem_0_4_W0_en = W0_en & _GEN_24;
  assign mem_0_4_W0_mask = W0_mask[4];
  assign mem_0_4_R0_addr = R0_addr[25:0];
  assign mem_0_4_R0_clk = R0_clk;
  assign _GEN_33 = R0_addr_sel == 2'h0;
  assign mem_0_4_R0_en = R0_en & _GEN_25;
  assign mem_0_5_W0_addr = W0_addr[25:0];
  assign mem_0_5_W0_clk = W0_clk;
  assign mem_0_5_W0_data = W0_data[47:40];
  assign _GEN_34 = W0_addr_sel == 2'h0;
  assign mem_0_5_W0_en = W0_en & _GEN_24;
  assign mem_0_5_W0_mask = W0_mask[5];
  assign mem_0_5_R0_addr = R0_addr[25:0];
  assign mem_0_5_R0_clk = R0_clk;
  assign _GEN_35 = R0_addr_sel == 2'h0;
  assign mem_0_5_R0_en = R0_en & _GEN_25;
  assign mem_0_6_W0_addr = W0_addr[25:0];
  assign mem_0_6_W0_clk = W0_clk;
  assign mem_0_6_W0_data = W0_data[55:48];
  assign _GEN_36 = W0_addr_sel == 2'h0;
  assign mem_0_6_W0_en = W0_en & _GEN_24;
  assign mem_0_6_W0_mask = W0_mask[6];
  assign mem_0_6_R0_addr = R0_addr[25:0];
  assign mem_0_6_R0_clk = R0_clk;
  assign _GEN_37 = R0_addr_sel == 2'h0;
  assign mem_0_6_R0_en = R0_en & _GEN_25;
  assign mem_0_7_W0_addr = W0_addr[25:0];
  assign mem_0_7_W0_clk = W0_clk;
  assign mem_0_7_W0_data = W0_data[63:56];
  assign _GEN_38 = W0_addr_sel == 2'h0;
  assign mem_0_7_W0_en = W0_en & _GEN_24;
  assign mem_0_7_W0_mask = W0_mask[7];
  assign mem_0_7_R0_addr = R0_addr[25:0];
  assign mem_0_7_R0_clk = R0_clk;
  assign _GEN_39 = R0_addr_sel == 2'h0;
  assign mem_0_7_R0_en = R0_en & _GEN_25;
  assign mem_1_0_W0_addr = W0_addr[25:0];
  assign mem_1_0_W0_clk = W0_clk;
  assign mem_1_0_W0_data = W0_data[7:0];
  assign _GEN_40 = W0_addr_sel == 2'h1;
  assign mem_1_0_W0_en = W0_en & _GEN_40;
  assign mem_1_0_W0_mask = W0_mask[0];
  assign mem_1_0_R0_addr = R0_addr[25:0];
  assign mem_1_0_R0_clk = R0_clk;
  assign _GEN_41 = R0_addr_sel == 2'h1;
  assign mem_1_0_R0_en = R0_en & _GEN_41;
  assign mem_1_1_W0_addr = W0_addr[25:0];
  assign mem_1_1_W0_clk = W0_clk;
  assign mem_1_1_W0_data = W0_data[15:8];
  assign _GEN_42 = W0_addr_sel == 2'h1;
  assign mem_1_1_W0_en = W0_en & _GEN_40;
  assign mem_1_1_W0_mask = W0_mask[1];
  assign mem_1_1_R0_addr = R0_addr[25:0];
  assign mem_1_1_R0_clk = R0_clk;
  assign _GEN_43 = R0_addr_sel == 2'h1;
  assign mem_1_1_R0_en = R0_en & _GEN_41;
  assign mem_1_2_W0_addr = W0_addr[25:0];
  assign mem_1_2_W0_clk = W0_clk;
  assign mem_1_2_W0_data = W0_data[23:16];
  assign _GEN_44 = W0_addr_sel == 2'h1;
  assign mem_1_2_W0_en = W0_en & _GEN_40;
  assign mem_1_2_W0_mask = W0_mask[2];
  assign mem_1_2_R0_addr = R0_addr[25:0];
  assign mem_1_2_R0_clk = R0_clk;
  assign _GEN_45 = R0_addr_sel == 2'h1;
  assign mem_1_2_R0_en = R0_en & _GEN_41;
  assign mem_1_3_W0_addr = W0_addr[25:0];
  assign mem_1_3_W0_clk = W0_clk;
  assign mem_1_3_W0_data = W0_data[31:24];
  assign _GEN_46 = W0_addr_sel == 2'h1;
  assign mem_1_3_W0_en = W0_en & _GEN_40;
  assign mem_1_3_W0_mask = W0_mask[3];
  assign mem_1_3_R0_addr = R0_addr[25:0];
  assign mem_1_3_R0_clk = R0_clk;
  assign _GEN_47 = R0_addr_sel == 2'h1;
  assign mem_1_3_R0_en = R0_en & _GEN_41;
  assign mem_1_4_W0_addr = W0_addr[25:0];
  assign mem_1_4_W0_clk = W0_clk;
  assign mem_1_4_W0_data = W0_data[39:32];
  assign _GEN_48 = W0_addr_sel == 2'h1;
  assign mem_1_4_W0_en = W0_en & _GEN_40;
  assign mem_1_4_W0_mask = W0_mask[4];
  assign mem_1_4_R0_addr = R0_addr[25:0];
  assign mem_1_4_R0_clk = R0_clk;
  assign _GEN_49 = R0_addr_sel == 2'h1;
  assign mem_1_4_R0_en = R0_en & _GEN_41;
  assign mem_1_5_W0_addr = W0_addr[25:0];
  assign mem_1_5_W0_clk = W0_clk;
  assign mem_1_5_W0_data = W0_data[47:40];
  assign _GEN_50 = W0_addr_sel == 2'h1;
  assign mem_1_5_W0_en = W0_en & _GEN_40;
  assign mem_1_5_W0_mask = W0_mask[5];
  assign mem_1_5_R0_addr = R0_addr[25:0];
  assign mem_1_5_R0_clk = R0_clk;
  assign _GEN_51 = R0_addr_sel == 2'h1;
  assign mem_1_5_R0_en = R0_en & _GEN_41;
  assign mem_1_6_W0_addr = W0_addr[25:0];
  assign mem_1_6_W0_clk = W0_clk;
  assign mem_1_6_W0_data = W0_data[55:48];
  assign _GEN_52 = W0_addr_sel == 2'h1;
  assign mem_1_6_W0_en = W0_en & _GEN_40;
  assign mem_1_6_W0_mask = W0_mask[6];
  assign mem_1_6_R0_addr = R0_addr[25:0];
  assign mem_1_6_R0_clk = R0_clk;
  assign _GEN_53 = R0_addr_sel == 2'h1;
  assign mem_1_6_R0_en = R0_en & _GEN_41;
  assign mem_1_7_W0_addr = W0_addr[25:0];
  assign mem_1_7_W0_clk = W0_clk;
  assign mem_1_7_W0_data = W0_data[63:56];
  assign _GEN_54 = W0_addr_sel == 2'h1;
  assign mem_1_7_W0_en = W0_en & _GEN_40;
  assign mem_1_7_W0_mask = W0_mask[7];
  assign mem_1_7_R0_addr = R0_addr[25:0];
  assign mem_1_7_R0_clk = R0_clk;
  assign _GEN_55 = R0_addr_sel == 2'h1;
  assign mem_1_7_R0_en = R0_en & _GEN_41;
  assign mem_2_0_W0_addr = W0_addr[25:0];
  assign mem_2_0_W0_clk = W0_clk;
  assign mem_2_0_W0_data = W0_data[7:0];
  assign _GEN_56 = W0_addr_sel == 2'h2;
  assign mem_2_0_W0_en = W0_en & _GEN_56;
  assign mem_2_0_W0_mask = W0_mask[0];
  assign mem_2_0_R0_addr = R0_addr[25:0];
  assign mem_2_0_R0_clk = R0_clk;
  assign _GEN_57 = R0_addr_sel == 2'h2;
  assign mem_2_0_R0_en = R0_en & _GEN_57;
  assign mem_2_1_W0_addr = W0_addr[25:0];
  assign mem_2_1_W0_clk = W0_clk;
  assign mem_2_1_W0_data = W0_data[15:8];
  assign _GEN_58 = W0_addr_sel == 2'h2;
  assign mem_2_1_W0_en = W0_en & _GEN_56;
  assign mem_2_1_W0_mask = W0_mask[1];
  assign mem_2_1_R0_addr = R0_addr[25:0];
  assign mem_2_1_R0_clk = R0_clk;
  assign _GEN_59 = R0_addr_sel == 2'h2;
  assign mem_2_1_R0_en = R0_en & _GEN_57;
  assign mem_2_2_W0_addr = W0_addr[25:0];
  assign mem_2_2_W0_clk = W0_clk;
  assign mem_2_2_W0_data = W0_data[23:16];
  assign _GEN_60 = W0_addr_sel == 2'h2;
  assign mem_2_2_W0_en = W0_en & _GEN_56;
  assign mem_2_2_W0_mask = W0_mask[2];
  assign mem_2_2_R0_addr = R0_addr[25:0];
  assign mem_2_2_R0_clk = R0_clk;
  assign _GEN_61 = R0_addr_sel == 2'h2;
  assign mem_2_2_R0_en = R0_en & _GEN_57;
  assign mem_2_3_W0_addr = W0_addr[25:0];
  assign mem_2_3_W0_clk = W0_clk;
  assign mem_2_3_W0_data = W0_data[31:24];
  assign _GEN_62 = W0_addr_sel == 2'h2;
  assign mem_2_3_W0_en = W0_en & _GEN_56;
  assign mem_2_3_W0_mask = W0_mask[3];
  assign mem_2_3_R0_addr = R0_addr[25:0];
  assign mem_2_3_R0_clk = R0_clk;
  assign _GEN_63 = R0_addr_sel == 2'h2;
  assign mem_2_3_R0_en = R0_en & _GEN_57;
  assign mem_2_4_W0_addr = W0_addr[25:0];
  assign mem_2_4_W0_clk = W0_clk;
  assign mem_2_4_W0_data = W0_data[39:32];
  assign _GEN_64 = W0_addr_sel == 2'h2;
  assign mem_2_4_W0_en = W0_en & _GEN_56;
  assign mem_2_4_W0_mask = W0_mask[4];
  assign mem_2_4_R0_addr = R0_addr[25:0];
  assign mem_2_4_R0_clk = R0_clk;
  assign _GEN_65 = R0_addr_sel == 2'h2;
  assign mem_2_4_R0_en = R0_en & _GEN_57;
  assign mem_2_5_W0_addr = W0_addr[25:0];
  assign mem_2_5_W0_clk = W0_clk;
  assign mem_2_5_W0_data = W0_data[47:40];
  assign _GEN_66 = W0_addr_sel == 2'h2;
  assign mem_2_5_W0_en = W0_en & _GEN_56;
  assign mem_2_5_W0_mask = W0_mask[5];
  assign mem_2_5_R0_addr = R0_addr[25:0];
  assign mem_2_5_R0_clk = R0_clk;
  assign _GEN_67 = R0_addr_sel == 2'h2;
  assign mem_2_5_R0_en = R0_en & _GEN_57;
  assign mem_2_6_W0_addr = W0_addr[25:0];
  assign mem_2_6_W0_clk = W0_clk;
  assign mem_2_6_W0_data = W0_data[55:48];
  assign _GEN_68 = W0_addr_sel == 2'h2;
  assign mem_2_6_W0_en = W0_en & _GEN_56;
  assign mem_2_6_W0_mask = W0_mask[6];
  assign mem_2_6_R0_addr = R0_addr[25:0];
  assign mem_2_6_R0_clk = R0_clk;
  assign _GEN_69 = R0_addr_sel == 2'h2;
  assign mem_2_6_R0_en = R0_en & _GEN_57;
  assign mem_2_7_W0_addr = W0_addr[25:0];
  assign mem_2_7_W0_clk = W0_clk;
  assign mem_2_7_W0_data = W0_data[63:56];
  assign _GEN_70 = W0_addr_sel == 2'h2;
  assign mem_2_7_W0_en = W0_en & _GEN_56;
  assign mem_2_7_W0_mask = W0_mask[7];
  assign mem_2_7_R0_addr = R0_addr[25:0];
  assign mem_2_7_R0_clk = R0_clk;
  assign _GEN_71 = R0_addr_sel == 2'h2;
  assign mem_2_7_R0_en = R0_en & _GEN_57;
  assign mem_3_0_W0_addr = W0_addr[25:0];
  assign mem_3_0_W0_clk = W0_clk;
  assign mem_3_0_W0_data = W0_data[7:0];
  assign _GEN_72 = W0_addr_sel == 2'h3;
  assign mem_3_0_W0_en = W0_en & _GEN_72;
  assign mem_3_0_W0_mask = W0_mask[0];
  assign mem_3_0_R0_addr = R0_addr[25:0];
  assign mem_3_0_R0_clk = R0_clk;
  assign _GEN_73 = R0_addr_sel == 2'h3;
  assign mem_3_0_R0_en = R0_en & _GEN_73;
  assign mem_3_1_W0_addr = W0_addr[25:0];
  assign mem_3_1_W0_clk = W0_clk;
  assign mem_3_1_W0_data = W0_data[15:8];
  assign _GEN_74 = W0_addr_sel == 2'h3;
  assign mem_3_1_W0_en = W0_en & _GEN_72;
  assign mem_3_1_W0_mask = W0_mask[1];
  assign mem_3_1_R0_addr = R0_addr[25:0];
  assign mem_3_1_R0_clk = R0_clk;
  assign _GEN_75 = R0_addr_sel == 2'h3;
  assign mem_3_1_R0_en = R0_en & _GEN_73;
  assign mem_3_2_W0_addr = W0_addr[25:0];
  assign mem_3_2_W0_clk = W0_clk;
  assign mem_3_2_W0_data = W0_data[23:16];
  assign _GEN_76 = W0_addr_sel == 2'h3;
  assign mem_3_2_W0_en = W0_en & _GEN_72;
  assign mem_3_2_W0_mask = W0_mask[2];
  assign mem_3_2_R0_addr = R0_addr[25:0];
  assign mem_3_2_R0_clk = R0_clk;
  assign _GEN_77 = R0_addr_sel == 2'h3;
  assign mem_3_2_R0_en = R0_en & _GEN_73;
  assign mem_3_3_W0_addr = W0_addr[25:0];
  assign mem_3_3_W0_clk = W0_clk;
  assign mem_3_3_W0_data = W0_data[31:24];
  assign _GEN_78 = W0_addr_sel == 2'h3;
  assign mem_3_3_W0_en = W0_en & _GEN_72;
  assign mem_3_3_W0_mask = W0_mask[3];
  assign mem_3_3_R0_addr = R0_addr[25:0];
  assign mem_3_3_R0_clk = R0_clk;
  assign _GEN_79 = R0_addr_sel == 2'h3;
  assign mem_3_3_R0_en = R0_en & _GEN_73;
  assign mem_3_4_W0_addr = W0_addr[25:0];
  assign mem_3_4_W0_clk = W0_clk;
  assign mem_3_4_W0_data = W0_data[39:32];
  assign _GEN_80 = W0_addr_sel == 2'h3;
  assign mem_3_4_W0_en = W0_en & _GEN_72;
  assign mem_3_4_W0_mask = W0_mask[4];
  assign mem_3_4_R0_addr = R0_addr[25:0];
  assign mem_3_4_R0_clk = R0_clk;
  assign _GEN_81 = R0_addr_sel == 2'h3;
  assign mem_3_4_R0_en = R0_en & _GEN_73;
  assign mem_3_5_W0_addr = W0_addr[25:0];
  assign mem_3_5_W0_clk = W0_clk;
  assign mem_3_5_W0_data = W0_data[47:40];
  assign _GEN_82 = W0_addr_sel == 2'h3;
  assign mem_3_5_W0_en = W0_en & _GEN_72;
  assign mem_3_5_W0_mask = W0_mask[5];
  assign mem_3_5_R0_addr = R0_addr[25:0];
  assign mem_3_5_R0_clk = R0_clk;
  assign _GEN_83 = R0_addr_sel == 2'h3;
  assign mem_3_5_R0_en = R0_en & _GEN_73;
  assign mem_3_6_W0_addr = W0_addr[25:0];
  assign mem_3_6_W0_clk = W0_clk;
  assign mem_3_6_W0_data = W0_data[55:48];
  assign _GEN_84 = W0_addr_sel == 2'h3;
  assign mem_3_6_W0_en = W0_en & _GEN_72;
  assign mem_3_6_W0_mask = W0_mask[6];
  assign mem_3_6_R0_addr = R0_addr[25:0];
  assign mem_3_6_R0_clk = R0_clk;
  assign _GEN_85 = R0_addr_sel == 2'h3;
  assign mem_3_6_R0_en = R0_en & _GEN_73;
  assign mem_3_7_W0_addr = W0_addr[25:0];
  assign mem_3_7_W0_clk = W0_clk;
  assign mem_3_7_W0_data = W0_data[63:56];
  assign _GEN_86 = W0_addr_sel == 2'h3;
  assign mem_3_7_W0_en = W0_en & _GEN_72;
  assign mem_3_7_W0_mask = W0_mask[7];
  assign mem_3_7_R0_addr = R0_addr[25:0];
  assign mem_3_7_R0_clk = R0_clk;
  assign _GEN_87 = R0_addr_sel == 2'h3;
  assign mem_3_7_R0_en = R0_en & _GEN_73;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  R0_addr_sel_reg = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge R0_clk) begin
    if (R0_en) begin
      R0_addr_sel_reg <= R0_addr_sel;
    end
  end
endmodule
module split_mem_ext(
  input  [25:0] W0_addr,
  input         W0_clk,
  input  [7:0]  W0_data,
  input         W0_en,
  input         W0_mask,
  input  [25:0] R0_addr,
  input         R0_clk,
  output [7:0]  R0_data,
  input         R0_en
);
  reg [7:0] ram [0:67108863];
  reg [31:0] _RAND_0;
  wire [7:0] ram_R_0_data;
  wire [25:0] ram_R_0_addr;
  wire [7:0] ram_W_0_data;
  wire [25:0] ram_W_0_addr;
  wire  ram_W_0_mask;
  wire  ram_W_0_en;
  wire  _GEN_0;
  wire [25:0] _GEN_1;
  reg [25:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_1;
  wire  ram_R_0_addr_en;
  wire  _GEN_2;
  wire  _GEN_3;
  wire [25:0] _GEN_4;
  wire [7:0] _GEN_5;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr];
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data;
  assign _GEN_0 = R0_en;
  assign _GEN_1 = R0_addr;
  assign ram_R_0_addr_en = R0_en;
  assign _GEN_2 = W0_en;
  assign _GEN_3 = W0_mask;
  assign _GEN_4 = W0_addr;
  assign _GEN_5 = W0_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 67108864; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_1[25:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data;
    end
  end
  always @(posedge R0_clk) begin
    if (_GEN_0) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule

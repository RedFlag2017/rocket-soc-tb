`include "../svtb/test/base_test.sv"
`include "../svtb/test/test_sanity01.sv"
`include "../svtb/test/test_demo.sv"



